// Global parameters

// ICA PARAMS
parameter DIMENSION = 5;
parameter SAMPLES = 1024;

// CORDIC CONSTS
parameter DATA_WIDTH = 32;
parameter CORDIC_WIDTH = 38;
parameter CORDIC_STAGES = 16;
parameter ANGLE_WIDTH = 16;