`timescale 1ns / 1ps

module tb_updateTop();

    parameter N = 5;
    parameter M = 8;
    parameter DATA_WIDTH = 32;
    parameter FRAC_WIDTH = 20;
    parameter CORDIC_WIDTH = 38;
    parameter ANGLE_WIDTH = 16;
    parameter CORDIC_STAGES = 16;
    parameter CLK_PERIOD = 10;
    parameter LOGM = 3;
    parameter ADDR_WIDTH = 10;

    reg clk;
    reg rst_n;
    reg nreset;
    reg en;
    reg [N*DATA_WIDTH-1:0] W_in;
    reg [N*M*DATA_WIDTH-1:0] Z_in;
    reg [1:0] scica_stage_in;
    
    // Z memory interface signals
    wire Z_in_en;
    wire [ADDR_WIDTH-1:0] Z_address1;
    wire [ADDR_WIDTH-1:0] Z_address2;
    wire signed [DATA_WIDTH-1:0] Z_in1;
    wire signed [DATA_WIDTH-1:0] Z_in2;
    wire Z_in_valid;
    reg zmem_writeEn;
    reg [ADDR_WIDTH-1:0] zmem_write_addr1;
    reg [ADDR_WIDTH-1:0] zmem_write_addr2;
    reg signed [DATA_WIDTH-1:0] zmem_din1;
    
    wire ica_cordic_vec_en;
    wire signed [DATA_WIDTH-1:0] ica_cordic_vec_xin;
    wire signed [DATA_WIDTH-1:0] ica_cordic_vec_yin;
    wire ica_cordic_vec_angle_calc_en;
    wire ica_cordic_rot1_en;
    wire signed [DATA_WIDTH-1:0] ica_cordic_rot1_xin;
    wire signed [DATA_WIDTH-1:0] ica_cordic_rot1_yin;
    wire signed [ANGLE_WIDTH-1:0] ica_cordic_rot1_angle_in;
    wire ica_cordic_rot1_angle_microRot_n;
    wire [CORDIC_STAGES-1:0] ica_cordic_rot1_microRot_ext_in;
    wire ica_cordic_rot1_microRot_ext_vld;
    wire [1:0] ica_cordic_rot1_quad_in;
    
    wire cordic_vec_opvld;
    wire signed [DATA_WIDTH-1:0] cordic_vec_xout;
    wire [1:0] cordic_vec_quad_out;
    wire cordic_vec_microRot_out_start;
    wire cordic_rot1_opvld;
    wire signed [DATA_WIDTH-1:0] cordic_rot1_xout;
    
    // Keep unused CORDIC outputs for the CORDIC wrapper
    wire [CORDIC_STAGES-1:0] cordic_vec_microRot_out;
    wire signed [ANGLE_WIDTH-1:0] cordic_vec_angle_out;
    wire signed [DATA_WIDTH-1:0] cordic_rot1_yout;
    wire cordic_rot2_opvld;
    wire signed [DATA_WIDTH-1:0] cordic_rot2_xout;
    wire signed [DATA_WIDTH-1:0] cordic_rot2_yout;
    wire ica_cordic_rot2_en;
    wire signed [DATA_WIDTH-1:0] ica_cordic_rot2_xin;
    wire signed [DATA_WIDTH-1:0] ica_cordic_rot2_yin;
    wire [1:0] ica_cordic_rot2_quad_in;
    wire [CORDIC_STAGES-1:0] ica_cordic_rot2_microRot_in;
    
    wire [N*DATA_WIDTH-1:0] W_out;
    wire output_valid;

    // Memory arrays to store test vectors
    reg [DATA_WIDTH-1:0] W_test [0:N-1];
    reg [DATA_WIDTH-1:0] Z_test [0:(N*M)-1];
    reg [DATA_WIDTH-1:0] expected [0:N-1];
    integer vector_count;
    integer i, j; // Loop variables
    
    // File handle for output
    integer output_file;

    initial begin
        clk = 0;
        forever #(CLK_PERIOD/2) clk = ~clk;
    end

    initial begin
        // Read the memory files generated by the Python script
        $readmemh("_W_in.mem", W_test);
        $readmemh("_Z_in.mem", Z_test);
        $readmemh("_expected.mem", expected);
        
        $dumpfile("tb_updateTop.vcd");
        $dumpvars(0, tb_updateTop);
        
        vector_count = 0;
        rst_n = 0; nreset = 0; en = 0; W_in = 0; Z_in = 0; scica_stage_in = 2'b01;
        zmem_writeEn = 0; zmem_write_addr1 = 0; zmem_write_addr2 = 0; 
        zmem_din1 = 0;
        #30;
        rst_n = 1; nreset = 1;
        #25;

        // Load Z memory - inline implementation
        $display("Loading Z data into memory...");
        zmem_writeEn = 1;
        #10;
        for (i = 0; i < (N*M); i = i + 1) begin
            zmem_write_addr1 = i;
            zmem_write_addr2 = 0; 
            zmem_din1 = Z_test[i];
            @(posedge clk);
        end
        
        zmem_writeEn = 0;
        $display("Z data loading complete.");
        #20;
        
        // Run test - inline implementation
        for (i = 0; i < N; i = i + 1)
            W_in[i*DATA_WIDTH +: DATA_WIDTH] = W_test[i];
        
        // $display("Starting test with:");
        // $display("W_in: %h", W_in);
        
        en = 1;
        wait (output_valid == 1);
        en = 0;
        
        $display("Test Results:");
        for (i = 0; i < N; i = i + 1) begin
            $display("Vector %0d, W[%0d] = %08x (Expected = %08x)", 
                    vector_count, i, W_out[i*DATA_WIDTH +: DATA_WIDTH], expected[i]);
        end
        
        // Open file for appending and write compact results
        output_file = $fopen("test_results.txt", "a");
        if (output_file != 0) begin
            // $fwrite(output_file, "V%0d: ", vector_count);
            for (i = 0; i < N; i = i + 1) begin
                $fwrite(output_file, "%08x  %08x\n", W_out[i*DATA_WIDTH +: DATA_WIDTH], expected[i]);
            end
            // $fwrite(output_file, "\n");
            $fclose(output_file);
        end
        
        vector_count = vector_count + 1;
        
        #100;
        $finish;
    end

    // Z Memory instantiation
    zmem #(
        .DATA_WIDTH(DATA_WIDTH),
        .ADDR_WIDTH(ADDR_WIDTH),
        .LATENCY(1),
        .M(M),
        .N(N)
    ) zmem_inst (
        .clk(clk),
        .rst_n(rst_n),
        .readEn(Z_in_en),
        .writeEn(zmem_writeEn),
        .addr1(zmem_writeEn ? zmem_write_addr1 : Z_address1),
        .addr2(zmem_writeEn ? zmem_write_addr2 : Z_address2),
        .din1(zmem_din1),
        .dout1(Z_in1),
        .dout2(Z_in2),
        .dout_valid(Z_in_valid)
    );

    // Updated updateTop instantiation
    updateTop #(
        .N(N), .M(M), .DATA_WIDTH(DATA_WIDTH), .FRAC_WIDTH(FRAC_WIDTH),
        .CORDIC_WIDTH(CORDIC_WIDTH), .ANGLE_WIDTH(ANGLE_WIDTH), 
        .CORDIC_STAGES(CORDIC_STAGES), .LOGM(LOGM), .ADDR_WIDTH(ADDR_WIDTH)
    ) uut_updateTop (
        .clk(clk), 
        .rst_n(rst_n), 
        .en(en), 
        .W_in(W_in),  
        .Z_in1(Z_in1),
        .Z_in2(Z_in2),
        .Z_in_valid(Z_in_valid),
        .cordic_vec_opvld(cordic_vec_opvld), 
        .cordic_vec_xout(cordic_vec_xout),
        .cordic_vec_quad_out(cordic_vec_quad_out),
        .cordic_vec_microRot_out_start(cordic_vec_microRot_out_start), 
        .cordic_rot1_opvld(cordic_rot1_opvld), 
        .cordic_rot1_xout(cordic_rot1_xout), 
        .ica_cordic_vec_en(ica_cordic_vec_en), 
        .ica_cordic_vec_xin(ica_cordic_vec_xin),
        .ica_cordic_vec_yin(ica_cordic_vec_yin), 
        .ica_cordic_vec_angle_calc_en(ica_cordic_vec_angle_calc_en),
        .ica_cordic_rot1_en(ica_cordic_rot1_en), 
        .ica_cordic_rot1_xin(ica_cordic_rot1_xin),
        .ica_cordic_rot1_yin(ica_cordic_rot1_yin), 
        .ica_cordic_rot1_angle_in(ica_cordic_rot1_angle_in),
        .ica_cordic_rot1_angle_microRot_n(ica_cordic_rot1_angle_microRot_n),
        .ica_cordic_rot1_microRot_ext_in(ica_cordic_rot1_microRot_ext_in),
        .ica_cordic_rot1_microRot_ext_vld(ica_cordic_rot1_microRot_ext_vld),
        .ica_cordic_rot1_quad_in(ica_cordic_rot1_quad_in),
        .Z_in_en(Z_in_en),
        .Z_address1(Z_address1),
        .Z_address2(Z_address2),
        .W_out(W_out), 
        .output_valid(output_valid)
    );

    SCICA_CORDIC_wrapper #(
        .DATA_WIDTH(DATA_WIDTH), .CORDIC_STAGES(CORDIC_STAGES), 
        .CORDIC_WIDTH(CORDIC_WIDTH), .ANGLE_WIDTH(ANGLE_WIDTH)
    ) dut_cordic (
        .clk(clk), .nreset(nreset), .scica_stage_in(scica_stage_in),
        .ica_cordic_vec_en(ica_cordic_vec_en), .ica_cordic_vec_xin(ica_cordic_vec_xin),
        .ica_cordic_vec_yin(ica_cordic_vec_yin), .ica_cordic_vec_angle_calc_en(ica_cordic_vec_angle_calc_en),
        .ica_cordic_rot1_en(ica_cordic_rot1_en), .ica_cordic_rot1_xin(ica_cordic_rot1_xin),
        .ica_cordic_rot1_yin(ica_cordic_rot1_yin), .ica_cordic_rot1_angle_in(ica_cordic_rot1_angle_in),
        .ica_cordic_rot1_angle_microRot_n(ica_cordic_rot1_angle_microRot_n),
        .ica_cordic_rot1_microRot_ext_in(ica_cordic_rot1_microRot_ext_in),
        .ica_cordic_rot1_microRot_ext_vld(ica_cordic_rot1_microRot_ext_vld),
        .ica_cordic_rot1_quad_in(ica_cordic_rot1_quad_in), .ica_cordic_rot2_en(ica_cordic_rot2_en),
        .ica_cordic_rot2_xin(ica_cordic_rot2_xin), .ica_cordic_rot2_yin(ica_cordic_rot2_yin),
        .ica_cordic_rot2_quad_in(ica_cordic_rot2_quad_in), .ica_cordic_rot2_microRot_in(ica_cordic_rot2_microRot_in),
        .cordic_vec_opvld(cordic_vec_opvld), .cordic_vec_xout(cordic_vec_xout),
        .cordic_vec_microRot_out(cordic_vec_microRot_out), .cordic_vec_quad_out(cordic_vec_quad_out),
        .cordic_vec_microRot_out_start(cordic_vec_microRot_out_start), .cordic_vec_angle_out(cordic_vec_angle_out),
        .cordic_rot1_opvld(cordic_rot1_opvld), .cordic_rot1_xout(cordic_rot1_xout), .cordic_rot1_yout(cordic_rot1_yout),
        .cordic_rot2_opvld(cordic_rot2_opvld), .cordic_rot2_xout(cordic_rot2_xout), .cordic_rot2_yout(cordic_rot2_yout)
    );

endmodule